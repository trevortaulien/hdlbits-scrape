module top_module( 
    input [99:0] in,
    output [99:0] out
);
​
endmodule
​
